`ifndef DATA_OP
`define DATA_OP

`define STATE_FUNC	2'd0
`define STATE_UP	2'd1
`define STATE_LOW	2'd2

`define FUNCT_PORTA	8'd65
`define FUNCT_PORTB	8'd66
`define FUNCT_PORTC	8'd67
`define FUNCT_PORTD	8'd68
`define FUNCT_DUTYC	8'd69
`define FUNCT_SCLKS	8'd83
`define FUNCT_SCLKF	8'd70
`define FUNCT_NONE	8'd0

`endif